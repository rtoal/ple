module HelloWorld;
  initial
    $display("Hello, world!");
endmodule